module mem_matrix;
    reg[31:0] a [255:0];
    reg[31:0] w [255:0];
    reg[31:0] b [255:0];

    integer MATRIX_SIZE = 16;

    integer i;
    integer j;
    real proper_state;
    real correcting = (2**15 / 2);

    integer f;

    initial begin
        
        for (i = 0; i < (MATRIX_SIZE*MATRIX_SIZE); i = i + 1) begin
            a[i] = i % 10;
        end

        for (i = (MATRIX_SIZE*MATRIX_SIZE -1); i >= 0; i = i - 1) begin
            w[i] = i % 10;
        end

        for (i = 0; i < (MATRIX_SIZE*MATRIX_SIZE); i = i + 1) begin
            b[i] = 0;
        end

        $display("INPUT");
        $display("---------------------------");
        for (i = 0; i < MATRIX_SIZE; i = i + 1) begin
            for (j = 0; j < MATRIX_SIZE; j = j + 1) begin
                $write("%d ", a[i * MATRIX_SIZE + j]);
            end
            $write("\n");
        end
        $display("---------------------------");

        $display("WEIGHTS");
        $display("---------------------------");
        for (i = 0; i < MATRIX_SIZE; i = i + 1) begin
            for (j = 0; j < MATRIX_SIZE; j = j + 1) begin
                $write("%d ", w[i * MATRIX_SIZE + j]);
            end
            $write("\n");
        end
        $display("---------------------------");

        $crossbar(16, a[0], a[1], a[2], a[3],
                    a[4], a[5], a[6], a[7],
                    a[8], a[9], a[10], a[11],
                    a[12], a[13], a[14], a[15], 
                    a[16], a[17], a[18], a[19],
                    a[20], a[21], a[22], a[23],
                    a[24], a[25], a[26], a[27],
                    a[28], a[29], a[30], a[31], 
                    a[32], a[33], a[34], a[35],
                    a[36], a[37], a[38], a[39],
                    a[40], a[41], a[42], a[43],
                    a[44], a[45], a[46], a[47], 
                    a[48], a[49], a[50], a[51],
                    a[52], a[53], a[54], a[55],
                    a[56], a[57], a[58], a[59],
                    a[60], a[61], a[62], a[63],
                    a[64], a[65], a[66], a[67],
                    a[68], a[69], a[70], a[71],
                    a[72], a[73], a[74], a[75],
                    a[76], a[77], a[78], a[79], 
                    a[80], a[81], a[82], a[83],
                    a[84], a[85], a[86], a[87],
                    a[88], a[89], a[90], a[91],
                    a[92], a[93], a[94], a[95], 
                    a[96], a[97], a[98], a[99],
                    a[100], a[101], a[102], a[103],
                    a[104], a[105], a[106], a[107],
                    a[108], a[109], a[110], a[111], 
                    a[112], a[113], a[114], a[115],
                    a[116], a[117], a[118], a[119],
                    a[120], a[121], a[122], a[123],
                    a[124], a[125], a[126], a[127],
                    a[128], a[129], a[130], a[131],
                    a[132], a[133], a[134], a[135],
                    a[136], a[137], a[138], a[139],
                    a[140], a[141], a[142], a[143], 
                    a[144], a[145], a[146], a[147],
                    a[148], a[149], a[150], a[151],
                    a[152], a[153], a[154], a[155],
                    a[156], a[157], a[158], a[159], 
                    a[160], a[161], a[162], a[163],
                    a[164], a[165], a[166], a[167],
                    a[168], a[169], a[170], a[171],
                    a[172], a[173], a[174], a[175], 
                    a[176], a[177], a[178], a[179],
                    a[180], a[181], a[182], a[183],
                    a[184], a[185], a[186], a[187],
                    a[188], a[189], a[190], a[191],
                    a[192], a[193], a[194], a[195],
                    a[196], a[197], a[198], a[199],
                    a[200], a[201], a[202], a[203],
                    a[204], a[205], a[206], a[207], 
                    a[208], a[209], a[210], a[211],
                    a[212], a[213], a[214], a[215],
                    a[216], a[217], a[218], a[219],
                    a[220], a[221], a[222], a[223], 
                    a[224], a[225], a[226], a[227],
                    a[228], a[229], a[230], a[231],
                    a[232], a[233], a[234], a[235],
                    a[236], a[237], a[238], a[239], 
                    a[240], a[241], a[242], a[243],
                    a[244], a[245], a[246], a[247],
                    a[248], a[249], a[250], a[251],
                    a[252], a[253], a[254], a[255],
                    w[0], w[1], w[2], w[3],
                    w[4], w[5], w[6], w[7],
                    w[8], w[9], w[10], w[11],
                    w[12], w[13], w[14], w[15], 
                    w[16], w[17], w[18], w[19],
                    w[20], w[21], w[22], w[23],
                    w[24], w[25], w[26], w[27],
                    w[28], w[29], w[30], w[31], 
                    w[32], w[33], w[34], w[35],
                    w[36], w[37], w[38], w[39],
                    w[40], w[41], w[42], w[43],
                    w[44], w[45], w[46], w[47], 
                    w[48], w[49], w[50], w[51],
                    w[52], w[53], w[54], w[55],
                    w[56], w[57], w[58], w[59],
                    w[60], w[61], w[62], w[63],
                    w[64], w[65], w[66], w[67],
                    w[68], w[69], w[70], w[71],
                    w[72], w[73], w[74], w[75],
                    w[76], w[77], w[78], w[79], 
                    w[80], w[81], w[82], w[83],
                    w[84], w[85], w[86], w[87],
                    w[88], w[89], w[90], w[91],
                    w[92], w[93], w[94], w[95], 
                    w[96], w[97], w[98], w[99],
                    w[100], w[101], w[102], w[103],
                    w[104], w[105], w[106], w[107],
                    w[108], w[109], w[110], w[111], 
                    w[112], w[113], w[114], w[115],
                    w[116], w[117], w[118], w[119],
                    w[120], w[121], w[122], w[123],
                    w[124], w[125], w[126], w[127],
                    w[128], w[129], w[130], w[131],
                    w[132], w[133], w[134], w[135],
                    w[136], w[137], w[138], w[139],
                    w[140], w[141], w[142], w[143], 
                    w[144], w[145], w[146], w[147],
                    w[148], w[149], w[150], w[151],
                    w[152], w[153], w[154], w[155],
                    w[156], w[157], w[158], w[159], 
                    w[160], w[161], w[162], w[163],
                    w[164], w[165], w[166], w[167],
                    w[168], w[169], w[170], w[171],
                    w[172], w[173], w[174], w[175], 
                    w[176], w[177], w[178], w[179],
                    w[180], w[181], w[182], w[183],
                    w[184], w[185], w[186], w[187],
                    w[188], w[189], w[190], w[191],
                    w[192], w[193], w[194], w[195],
                    w[196], w[197], w[198], w[199],
                    w[200], w[201], w[202], w[203],
                    w[204], w[205], w[206], w[207], 
                    w[208], w[209], w[210], w[211],
                    w[212], w[213], w[214], w[215],
                    w[216], w[217], w[218], w[219],
                    w[220], w[221], w[222], w[223], 
                    w[224], w[225], w[226], w[227],
                    w[228], w[229], w[230], w[231],
                    w[232], w[233], w[234], w[235],
                    w[236], w[237], w[238], w[239], 
                    w[240], w[241], w[242], w[243],
                    w[244], w[245], w[246], w[247],
                    w[248], w[249], w[250], w[251],
                    w[252], w[253], w[254], w[255],
                    b[0], b[1], b[2], b[3],
                    b[4], b[5], b[6], b[7],
                    b[8], b[9], b[10], b[11],
                    b[12], b[13], b[14], b[15], 
                    b[16], b[17], b[18], b[19],
                    b[20], b[21], b[22], b[23],
                    b[24], b[25], b[26], b[27],
                    b[28], b[29], b[30], b[31], 
                    b[32], b[33], b[34], b[35],
                    b[36], b[37], b[38], b[39],
                    b[40], b[41], b[42], b[43],
                    b[44], b[45], b[46], b[47], 
                    b[48], b[49], b[50], b[51],
                    b[52], b[53], b[54], b[55],
                    b[56], b[57], b[58], b[59],
                    b[60], b[61], b[62], b[63],
                    b[64], b[65], b[66], b[67],
                    b[68], b[69], b[70], b[71],
                    b[72], b[73], b[74], b[75],
                    b[76], b[77], b[78], b[79], 
                    b[80], b[81], b[82], b[83],
                    b[84], b[85], b[86], b[87],
                    b[88], b[89], b[90], b[91],
                    b[92], b[93], b[94], b[95], 
                    b[96], b[97], b[98], b[99],
                    b[100], b[101], b[102], b[103],
                    b[104], b[105], b[106], b[107],
                    b[108], b[109], b[110], b[111], 
                    b[112], b[113], b[114], b[115],
                    b[116], b[117], b[118], b[119],
                    b[120], b[121], b[122], b[123],
                    b[124], b[125], b[126], b[127],
                    b[128], b[129], b[130], b[131],
                    b[132], b[133], b[134], b[135],
                    b[136], b[137], b[138], b[139],
                    b[140], b[141], b[142], b[143], 
                    b[144], b[145], b[146], b[147],
                    b[148], b[149], b[150], b[151],
                    b[152], b[153], b[154], b[155],
                    b[156], b[157], b[158], b[159], 
                    b[160], b[161], b[162], b[163],
                    b[164], b[165], b[166], b[167],
                    b[168], b[169], b[170], b[171],
                    b[172], b[173], b[174], b[175], 
                    b[176], b[177], b[178], b[179],
                    b[180], b[181], b[182], b[183],
                    b[184], b[185], b[186], b[187],
                    b[188], b[189], b[190], b[191],
                    b[192], b[193], b[194], b[195],
                    b[196], b[197], b[198], b[199],
                    b[200], b[201], b[202], b[203],
                    b[204], b[205], b[206], b[207], 
                    b[208], b[209], b[210], b[211],
                    b[212], b[213], b[214], b[215],
                    b[216], b[217], b[218], b[219],
                    b[220], b[221], b[222], b[223], 
                    b[224], b[225], b[226], b[227],
                    b[228], b[229], b[230], b[231],
                    b[232], b[233], b[234], b[235],
                    b[236], b[237], b[238], b[239], 
                    b[240], b[241], b[242], b[243],
                    b[244], b[245], b[246], b[247],
                    b[248], b[249], b[250], b[251],
                    b[252], b[253], b[254], b[255]
                    );
        
        $display("OUTPUT");
        $display("---------------------------");
        for (i = 0; i < MATRIX_SIZE; i = i + 1) begin
            for (j = 0; j < MATRIX_SIZE; j = j + 1) begin
                $write("%d ", b[i * MATRIX_SIZE + j]);
            end
            $write("\n");
        end
        $display("---------------------------");
        
    end

endmodule