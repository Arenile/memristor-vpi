module mem_matrix;
    reg[31:0] a [63:0];
    reg[31:0] w [63:0];
    reg[31:0] b [63:0];

    integer MATRIX_SIZE = 8;

    integer i;
    integer j;
    real proper_state;
    real correcting = (2**15 / 2);

    integer f;

    initial begin
        a[0] = 9; a[1] = 2; a[2] = 2; a[3] = 5; a[4] = 3; a[5] = 6; a[6] = 6; a[7] = 8;
        a[8] = 2; a[9] = 1; a[10] = 9; a[11] = 2; a[12] = 8; a[13] = 5; a[14] = 6; a[15] = 5;
        a[16] = 9; a[17] = 2; a[18] = 2; a[19] = 5; a[20] = 3; a[21] = 6; a[22] = 6; a[23] = 8;
        a[24] = 2; a[25] = 1; a[26] = 9; a[27] = 2; a[28] = 8; a[29] = 5; a[30] = 6; a[31] = 5;
        a[32] = 9; a[33] = 2; a[34] = 2; a[35] = 5; a[36] = 3; a[37] = 6; a[38] = 6; a[39] = 8;
        a[40] = 2; a[41] = 1; a[42] = 9; a[43] = 2; a[44] = 8; a[45] = 5; a[46] = 6; a[47] = 5;
        a[48] = 9; a[49] = 2; a[50] = 2; a[51] = 5; a[52] = 3; a[53] = 6; a[54] = 6; a[55] = 8;
        a[56] = 2; a[57] = 1; a[58] = 9; a[59] = 2; a[60] = 8; a[61] = 5; a[62] = 6; a[63] = 5;

        w[0] = 6; w[1] = 3; w[2] = 2; w[3] = 3; w[4] = 8; w[5] = 3; w[6] = 5; w[7] = 1;
        w[8] = 2; w[9] = 1; w[10] = 5; w[11] = 2; w[12] = 8; w[13] = 5; w[14] = 6; w[15] = 5;
        w[16] = 5; w[17] = 3; w[18] = 2; w[19] = 5; w[20] = 3; w[21] = 6; w[22] = 4; w[23] = 8;
        w[24] = 7; w[25] = 2; w[26] = 8; w[27] = 7; w[28] = 8; w[29] = 5; w[30] = 6; w[31] = 2;
        w[32] = 8; w[33] = 4; w[34] = 2; w[35] = 1; w[36] = 3; w[37] = 3; w[38] = 3; w[39] = 5;
        w[40] = 1; w[41] = 1; w[42] = 9; w[43] = 6; w[44] = 8; w[45] = 5; w[46] = 4; w[47] = 4;
        w[48] = 1; w[49] = 2; w[50] = 3; w[51] = 3; w[52] = 3; w[53] = 5; w[54] = 8; w[55] = 8;
        w[56] = 2; w[57] = 1; w[58] = 3; w[59] = 4; w[60] = 8; w[61] = 5; w[62] = 9; w[63] = 5;

        for (i = 0; i < 16; i = i + 1) begin
            b[i] = 0;
        end

        $display("INPUT");
        $display("---------------------------");
        for (i = 0; i < MATRIX_SIZE; i = i + 1) begin
            for (j = 0; j < MATRIX_SIZE; j = j + 1) begin
                $write("%d ", a[i * MATRIX_SIZE + j]);
            end
            $write("\n");
        end
        $display("---------------------------");

        $display("WEIGHTS");
        $display("---------------------------");
        for (i = 0; i < MATRIX_SIZE; i = i + 1) begin
            for (j = 0; j < MATRIX_SIZE; j = j + 1) begin
                $write("%d ", w[i * MATRIX_SIZE + j]);
            end
            $write("\n");
        end
        $display("---------------------------");

        $crossbar(8, a[0], a[1], a[2], a[3],
                    a[4], a[5], a[6], a[7],
                    a[8], a[9], a[10], a[11],
                    a[12], a[13], a[14], a[15], 
                    a[16], a[17], a[18], a[19],
                    a[20], a[21], a[22], a[23],
                    a[24], a[25], a[26], a[27],
                    a[28], a[29], a[30], a[31], 
                    a[32], a[33], a[34], a[35],
                    a[36], a[37], a[38], a[39],
                    a[40], a[41], a[42], a[43],
                    a[44], a[45], a[46], a[47], 
                    a[48], a[49], a[50], a[51],
                    a[52], a[53], a[54], a[55],
                    a[56], a[57], a[58], a[59],
                    a[60], a[61], a[62], a[63],
                    w[0], w[1], w[2], w[3],
                    w[4], w[5], w[6], w[7],
                    w[8], w[9], w[10], w[11],
                    w[12], w[13], w[14], w[15], 
                    w[16], w[17], w[18], w[19],
                    w[20], w[21], w[22], w[23],
                    w[24], w[25], w[26], w[27],
                    w[28], w[29], w[30], w[31], 
                    w[32], w[33], w[34], w[35],
                    w[36], w[37], w[38], w[39],
                    w[40], w[41], w[42], w[43],
                    w[44], w[45], w[46], w[47], 
                    w[48], w[49], w[50], w[51],
                    w[52], w[53], w[54], w[55],
                    w[56], w[57], w[58], w[59],
                    w[60], w[61], w[62], w[63],
                    b[0], b[1], b[2], b[3],
                    b[4], b[5], b[6], b[7],
                    b[8], b[9], b[10], b[11],
                    b[12], b[13], b[14], b[15], 
                    b[16], b[17], b[18], b[19],
                    b[20], b[21], b[22], b[23],
                    b[24], b[25], b[26], b[27],
                    b[28], b[29], b[30], b[31], 
                    b[32], b[33], b[34], b[35],
                    b[36], b[37], b[38], b[39],
                    b[40], b[41], b[42], b[43],
                    b[44], b[45], b[46], b[47], 
                    b[48], b[49], b[50], b[51],
                    b[52], b[53], b[54], b[55],
                    b[56], b[57], b[58], b[59],
                    b[60], b[61], b[62], b[63]);
        
        $display("OUTPUT");
        $display("---------------------------");
        for (i = 0; i < MATRIX_SIZE; i = i + 1) begin
            for (j = 0; j < MATRIX_SIZE; j = j + 1) begin
                $write("%d ", b[i * MATRIX_SIZE + j]);
            end
            $write("\n");
        end
        $display("---------------------------");
        
    end

endmodule